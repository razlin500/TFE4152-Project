//-----------------------------------------------------------------------------
//
// Title       : getAlpha
// Design      : tsetlin
// Author      : 
// Company     : 
//
//-----------------------------------------------------------------------------
//
// File        : c:\My_Designs\TFE4152\tsetlin\src\getAlpha.v
// Generated   : Thu Oct 30 11:05:02 2025
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {getAlpha}}
module getAlpha ( b2 ,b1 ,b0 ,alpha );

output alpha ;
wire alpha ;

input b2 ;
wire b2 ;
input b1 ;
wire b1 ;
input b0 ;
wire b0 ;

//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule

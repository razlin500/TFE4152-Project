//-----------------------------------------------------------------------------
//
// Title       : register
// Design      : tsetlin
// Author      : 
// Company     : 
//
//-----------------------------------------------------------------------------
//
// File        : c:\My_Designs\TFE4152\tsetlin\src\register.v
// Generated   : Thu Oct 30 11:03:13 2025
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {register}}
module register ( b2 ,b1 ,b0 ,b2o ,b1o ,b0o ,clk );

output b2o ;
wire b2o ;
output b1o ;
wire b1o ;
output b0o ;
wire b0o ;

input b2 ;
wire b2 ;
input b1 ;
wire b1 ;
input b0 ;
wire b0 ;
input clk ;
wire clk ;

//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule

[aimspice]
[description]
364
*Current mirror
.include p18_cmos_models_tt.inc

.param length=0.5u width=4.63u 

Vdd 1 0 1.0V

Vout 6 0 1.0V


IB 1 2 45u

Iin 1 4 50u


M1 6 2 7 0 NMOS L=length W=width

M2 7 4 0 0 NMOS L=0.5length W=0.5width

M3 5 4 0 0 NMOS L=0.5length W=0.5width

M4 4 2 5 0 NMOS L=length W=width

M5 2 2 0 0 NMOS L=length W=0.25width

.plot dc id(M1)
[dc]
1
Vout
0
1
0.001
[ana]
1 0
[end]

[aimspice]
[description]
354
*Current mirror
.include p18_cmos_models_tt.inc

.param length=1u width=9.26u

Vdd 1 0 1.0V

Vout 6 0 1.0V



Ibias 1 2 45u

Iin 1 3 45u


M1 6 2 4 0 NMOS L=length W=0.25width

M2 4 3 0 0 NMOS L=length W=width

M3 5 3 0 0 NMOS L=length W=width

M4 3 2 5 0 NMOS L=length W=width

M5 2 2 0 0 NMOS L=length W=width

.plot dc id(M1)
[end]

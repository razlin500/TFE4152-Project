//-----------------------------------------------------------------------------
//
// Title       : D_flip_flop
// Design      : tsetlin
// Author      : Rasmus Nummelin
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : C:/Users/razli/ikke_onedrive/H2025/TFE4152/TFE4152-Project/Digital/tsetlin/src/D_flip_flop.v
// Generated   : Mon Nov  3 11:13:53 2025
// From        : Interface description file
// By          : ItfToHdl ver. 1.0
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps

//{{ Section below this comment is automatically maintained
//    and may be overwritten
//{module {D_flip_flop}}

module D_flip_flop ( D ,CLK ,Q ,Not_Q );

input D;
wire D;
input CLK;
wire CLK;
output Q;
wire Q;
output Not_Q;
wire Not_Q;

//}} End of automatically maintained section

// Enter your statements here //

endmodule

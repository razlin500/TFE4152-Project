[aimspice]
[description]
372
*Current mirror
.include p18_cmos_models_ff.inc

.param length=0.5u width=4.63u 

*Vdd 1 0 1.0V

Vout 6 0 1.0V


IB 1 2 dc 45u

Iin 1 4 50u


M1 6 2 7 0 NMOS L=length W=width

M2 7 4 0 0 NMOS L={length/2} W={width/2}

M3 5 4 0 0 NMOS L={length/2} W={width/2}

M4 4 2 5 0 NMOS L=length W=width

M5 2 2 0 0 NMOS L=length W={width/4}

.plot dc id(M1)
[options]
1
Tnom 50
[dc]
1
Iin
40u
50u
0.01u
[ana]
1 0
[end]

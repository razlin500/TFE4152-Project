[aimspice]
[description]
440
* Wide-swing cascode current

.include p18_cmos_models_tt.inc
.include p18_model_card.inc

.param length=1U
.param width=9.26U

Vdd1 3 0 dc 1.0V 
Vout 7 0 dc 1.0V

I_bias 3 1 dc 50u
I_in 3 2 dc 50u

MN1 7 5 6 0 NMOS L=length W=width
MN2 6 4 0 0 NMOS L=length W=width
MN3 8 2 0 4 NMOS L=length W=width
MN4 2 1 8 5 NMOS L=length W=width PD=500u PS=500u
MN5 1 1 0 0 NMOS L=length W=0.25width PD=500u PS=500u


.plot i(MN1)
[options]
1
Gmin 1.0E-38
[dc]
1
Vout
0
1
0.01
[ana]
1 1
0
1 1
1 1 0 5
1
i(vout)
[end]

[aimspice]
[description]
364
currentmirror
.param .param proc_delta = 0.95
vt_shift = 0.1
.include p18_model_card.inc
VDD vdd 0 2 DC
isrc Iin iin vdd


R1 vdd vx 122400
* DRAIN GATE BULK SOURCE
M1 M2 vx vx 0 out 0 NMOS W=5u L=1u
vx 0 0 NMOS W=5u L=1u
VOUT out 0 DC 0.9
*.op
.dc VOUT 0.5 1.5 0.01
.plot id(m2)
*.plot i(M2)
*.print i(M2)
.end

PHAT iin iin 0 0 NMOS 1/(n+1)^2
[end]

//-----------------------------------------------------------------------------
//
// Title       : combinatorics
// Design      : TsetlinMachine
// Author      : Rasmus Nummelin
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : C:/Users/razli/ikke_onedrive/H2025/TFE4152/TFE4152-Project/Digital/TsetlinMachine/TsetlinMachine/src/combinatorics.v
// Generated   : Mon Nov  3 12:23:53 2025
// From        : Interface description file
// By          : ItfToHdl ver. 1.0
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps

//{{ Section below this comment is automatically maintained
//    and may be overwritten
//{module {combinatorics}}

module combinatorics ( beta ,b0 ,b1 ,b2 ,b0o ,b1o ,b2o ,alpha );

input beta;
wire beta;
input b0;
wire b0;
input b1;
wire b1;
input b2;
wire b2;
output b0o;
wire b0o;
output b1o;
wire b1o;
output b2o;
wire b2o;
output alpha;
wire alpha;

//}} End of automatically maintained section

// Added some more text here

// Enter your statements here //

endmodule

//-----------------------------------------------------------------------------
//
// Title       : combinatorics
// Design      : tsetlin
// Author      : 
// Company     : 
//
//-----------------------------------------------------------------------------
//
// File        : c:\My_Designs\TFE4152\tsetlin\src\combinatorics.v
// Generated   : Thu Oct 30 10:59:53 2025
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {combinatorics}}
module combinatorics ( beta ,b2 ,b1 ,b0 ,b2o ,b1o ,b0o );

output b2o ;
wire b2o ;
output b1o ;
wire b1o ;
output b0o ;
wire b0o ;

input beta ;
wire beta ;
input b2 ;
wire b2 ;
input b1 ;
wire b1 ;
input b0 ;
wire b0 ;

//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule

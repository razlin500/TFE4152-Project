//-----------------------------------------------------------------------------
//
// Title       : Tsetlin_machine
// Design      : tsetlin
// Author      : NTNU
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : m:\TFE4152-Project\Digital\tsetlin\compile\Tsetlin machine.v
// Generated   : Mon Nov  3 10:52:51 2025
// From        : m:\TFE4152-Project\Digital\tsetlin\src\Tsetlin machine.bde
// By          : Bde2Verilog ver. 2.01
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`ifdef _VCP
`else
`define library(a,b)
`endif


// ---------- Design Unit Header ---------- //
`timescale 1ps / 1ps

module \\Tsetlin_machine (beta,alpha) ;

// ------------ Port declarations --------- //
input beta;
wire beta;
output alpha;
wire alpha;

endmodule 
